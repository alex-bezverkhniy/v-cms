module main

const (
	default_page_size = 10
	operations = {
		'neq': '!=', 
		'eq': '=', 
		'gt': '>', 
		'lt': '<', 
		'ge': '>=', 
		'le': '<=', 
		'like':'like', 
		'in':'in'
	}
)