module main

const (
	default_page_size = 10
)